module top_module( 
    input a,b, 
    output out );
    
    nor(out,a,b);

endmodule
