module top_module( 
    input a,b, 
    output out );
    
    and(out,a,b);

endmodule
