module top_module ( input x, y, output z );
    xnor(z,x,y);
endmodule
