module top_module( 
    input a,b, 
    output out );
    
    xnor(out,a,b);

endmodule
